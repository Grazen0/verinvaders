`ifndef INVADERS_NES_BRIDGE_VH
`define INVADERS_NES_BRIDGE_VH

`define JOYP_RIGHT 0
`define JOYP_LEFT 1
`define JOYP_DOWN 2
`define JOYP_UP 3
`define JOYP_START 4
`define JOYP_SELECT 5
`define JOYP_B 6
`define JOYP_A 7

`endif
